module moduleName (
    input wire [31:0] PC_adr
);
    
endmodule