module and (
    input wire A,
    input wire B,
    output wire Q
);

assign Q=A&B;

endmodule