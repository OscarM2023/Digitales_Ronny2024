`timescale 1ns/1ns
`include "signextend.sv"

module signextend_tb (
);
    reg [31:0] IN;
    wire [31:0] OUT;

signextend signextend_tb (

    .IN(IN),
    .OUT(OUT)
);
initial begin
    
    $dumpfile("signextend_tb.vcd");
    $dumpvars(0, signextend_tb);

    //lw
    IN = 32'b00000000000000000001000000000011;
    #10
    //OUT = 00000000_00000000_00000000_00000000

    IN = 32'b11111111111100000000000000000011; 
    #10;
    //OUT = 11111111_11111111_11111111_11111111


    //sw
    IN = 32'b00000000000000000001000000100011; 
    #10;
    //OUT = 00000000_00000000_00000000_00000000

    IN = 32'b11111110000000000001000000100011; 
    #10;
    //OUT = 11111111_11111111_11111111_11100000



    //beq
    IN = 32'b00000000000000000001000001100011; 
    #10;
    //OUT = 00000000_00000000_00000000_00000000

    IN = 32'b11111110000000000001000001100011; 
    #10;
    //OUT = 11111111_11111111_11111011_11110000



    //default
    IN = 32'b11111111111111111111111111111111; 
    #10;
    //OUT = 00000000_00000000_00000000_00000000

    $display("Test completado");
    $finish;



end




endmodule