module deco (
    ports
);
    
endmodule