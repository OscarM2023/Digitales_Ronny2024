module #(parameter WIDTH=32) (
    input wire [WIDTH-1:0] INSTRUCTION,

    output wire [3:0] ALUOP,
    output wire PCSRC, ALUSRC, MEMTOREAD, MEMWRITE, MEMTOREG, REGWRITE
);
    
//logica

endmodule