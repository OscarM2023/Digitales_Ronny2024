module hazard_unit (
    input wire MEMREAD_ID_EX,
    input wire [4:0] ARS1_IF_ID, ARS2_IF_ID, ARD_ID_EX,

    output wire STALL, MUX_SEL
);
    
//logica

endmodule